--Author: Mehran Goli
--Version: 1.0
--Date: 17-8-2019
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY reg_unit IS
                  
            PORT (regaddrs1,regaddrs2,writregaddrs : IN std_logic_vector(4 DOWNTO 0);
                  data_in : IN std_logic_vector(31 DOWNTO 0);
			      write_en,clk,clr : IN std_logic;
				  data_out1,data_out2 : OUT std_logic_vector(31 DOWNTO 0)
				  );
END;
ARCHITECTURE my_reg OF reg_unit IS
TYPE mymemory  IS ARRAY (0 TO 31) OF std_logic_vector(31 DOWNTO 0);
SIGNAL reg  :mymemory:=("00000000000000000000000000000001","00000000000000000000000000000111","00000000000000000000000000000011",
"00000000000000000000000000000001","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000");  
BEGIN
reg_p : PROCESS (clk,clr)
	    BEGIN
		    IF clr = '1' THEN
                reg <= (OTHERS =>( OTHERS => '0'));			
		    ELSIF clk'EVENT AND (clk = '1') AND( write_en = '1' )THEN
			    reg(conv_integer(writregaddrs)) <= data_in;
			END IF;	    
		END PROCESS reg_p;
		
--com_p : PROCESS (regaddrs1,regaddrs2)
	    --BEGIN
			  data_out1 <= reg(conv_integer(regaddrs1));
			  data_out2 <= reg(conv_integer(regaddrs2));   
		--END PROCESS com_p;		
END my_reg;

---------------------------------------------------------------
