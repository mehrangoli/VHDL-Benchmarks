--Author: Mehran Goli
--Version: 1.0
--Date: 17-8-2019
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY data_memory IS
    PORT (                 
                 address     : IN  std_logic_vector(4  DOWNTO 0);
                 data_in     : IN  std_logic_vector(31 DOWNTO 0);
                 mem_rw      : IN  std_logic;
                 clk, nrst   : IN  std_logic;       
                 data_out    : OUT std_logic_vector(31 DOWNTO 0)
         );
END data_memory;

ARCHITECTURE data_mem OF data_memory IS

     TYPE   memory IS ARRAY (0 TO 31) OF std_logic_vector(31 DOWNTO 0) ;          
     SIGNAL data_memory  :memory :=("00000000000000000000000000000011","00000000000000000000000000000001","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000");  
     
BEGIN
        PROCESS (clk,nrst)
        BEGIN
           -- IF nrst='0' THEN
                --data_memory <= (OTHERS => X"00000000");
            IF clk'EVENT AND clk='1' THEN
                IF mem_rw='1' THEN
                    data_out <= data_memory(conv_integer (address));
                ELSE
                    data_memory(conv_integer (address)) <= data_in;
                END IF;    
            END IF;
        END PROCESS;
END data_mem;   
