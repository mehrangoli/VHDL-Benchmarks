--Author: Mehran Goli
--Version: 1.0
--Date: 17-8-2019
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;

ENTITY instruction_memory IS
    PORT (
                 addr        : IN  std_logic_vector(4  DOWNTO 0);
                 clk, nrst   : IN  std_logic;   
                 instr       : OUT std_logic_vector(31 DOWNTO 0)                
         );
END instruction_memory;

ARCHITECTURE instr_mem OF instruction_memory IS

     TYPE   memory IS ARRAY (0 TO 31) OF std_logic_vector(31 DOWNTO 0) ;          
     SIGNAL instr_memory  :memory :=("00000000000000010001000000100000","00000000000000010001100000100001","00000000000000010010000000100010",
     "00000000000000010010100000100011","00000000000000010011000000100100","00000000000000010011100000100101","00000000000000010100000000100110",
     "00000000000000010100100000101010","00000000000000010101000000101011","00000000000000010101100000000110","00000000000000010110000000000100",
     "00000000000000010110100000001000","00100000000011100000000000000001","00100100000100010000000000000010","00110000000100100000000000000111",
     "00010000000100110000000000000001","00010100000101000000000000000001","00001000000101010000000000000010","10000000000101100000000000000010",
     "10001100000110000000000000000001","00110100000110010000000000000111","10100000000110100000000000000001","00101000000110110000000000000010",
     "00101100000111000000000000001011","10101100000111010000000000000001","00111000000111110000000000000111","00000000000000000000000000000000",
     "00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000","00000000000000000000000000000000",
     "00000000000000000000000000000000");  
     
BEGIN
        PROCESS (clk)
        BEGIN
           -- IF nrst='0' THEN
              --  instr_memory <= (OTHERS => X"00000000");
            IF clk'EVENT AND clk='1' THEN
                instr <= instr_memory(conv_integer (addr));
            END IF;
        END PROCESS;
END instr_mem;        
